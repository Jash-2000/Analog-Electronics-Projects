
.model BC108A NPN(Is=7.049f Xti=3 Eg=1.11 Vaf=116.3 Bf=375.5 Ise=7.049f Ne=1.281 Ikf=4.589 Nk=.5 Xtb=1.5 Br=2.611 Isc=121.7p Nc=1.865 Ikr=5.313 Rc=1.464 Cjc=5.38p Mjc=.329 Vjc=.6218 Fc=.5 Cje=11.5p Mje=.2717 Vje=.5 Tr=10n Tf=451p Itf=6.194 Xtf=17.43 Vtf=10)

RC 1 2 20K
R3 3 0 50K
RE 4 5 1K
CL 2 0 10N
Q1 2 3 4 BC108A
VCB 1 0 10
VEB1 5 6 -1
VEB 6 0 sin(0 10m 1K)AC

.op
.DC VEB
.AC DEC 50 10 10Meg
.step Param x -1.6 -0.4 0.12
.tran 0.02 5m
.END
